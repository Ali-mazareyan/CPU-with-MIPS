
module MEM_Dastoorat(Reset,AR,OUT);
input Reset;
input [15:0] AR;
output reg [31:0] OUT;

reg [15:0] H [0:65535];
integer i;

always @(*)
begin
	if(Reset==1)
	begin
		OUT = 0;
		H[0]=16'b0000010011101000; 
		H[1]=16'b0000000000000001; 
		//Add AC,1256	
		H[2]=16'b0000001100100000;
		H[3]=16'b0000000000000010;
		//Sub AC,800
		H[4]=16'b0001101110001101;
		H[5]=16'b0000000000000100;
		//AND AC,7053
		H[6]=16'b0000000011111111;
		H[7]=16'b0000000000001000;
		//OR AC,255
		H[8]=16'b0010101011110001;
		H[9]=16'b0000000000010000;
		//XOR AC,10993
		H[10]=16'b0000000000000011;
		H[11]=16'b0000000000100000;
		//AC , Shift Rast (3 Bit)
		H[12]=16'b0000000000000010;
		H[13]=16'b0000000001000000;
		//AC , Shift Chap (2Bit)
		H[14]=16'b0000000000000000;
		H[15]=16'b0000000010000000;
		//AC , NOT	
		H[16]=16'b0000000000001001;
		H[17]=16'b0000000100000000;		
		//Write AC,CH[9]
		H[18]=16'b0000000000001001;
		H[19]=16'b0000001000000000;	
		//Print(OR),CH[9]

		for (i=20;i<65536;i=i+1)
			H[i]=16'b0;		
	end
	else
	begin
		OUT = {H[AR+1],H[AR]};
	end


end


endmodule
